module addition(input [23:0] a, output [23:0] done);
    assign done = a + 2;
endmodule
